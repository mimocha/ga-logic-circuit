// Input != Output

module flip (
	input wire IN,
	output wire OUT
	);
	
//	OUT != IN;
	
endmodule 
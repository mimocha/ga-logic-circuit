// Input == Output

module linear (
	input wire IN,
	input wire A,
	output wire OUT
	);
	
assign	OUT = IN;
	
endmodule 
// fpga_main.v

module fpga_main (
	input	IN,
	output	OUT
	);
	
	assign OUT = IN;

endmodule 
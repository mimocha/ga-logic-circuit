// Input == Output

module linear (
	input wire IN,
	output wire OUT
	);
	
assign	OUT = IN;
	
endmodule 
/*--------------------------------------------------------------------------//
// Original Title:        de0_nano_soc_baseline.v                           //
// Rev:                   Rev 0.1                                           //
// Last Revised:          09/14/2015                                        //
//--------------------------------------------------------------------------//
// Description: Baseline design file contains DE0 Nano SoC                  //
//              Board pins and I/O Standards.                               //
//--------------------------------------------------------------------------//
//Copyright 2015 Altera Corporation. All rights reserved.  Altera products
//are protected under numerous U.S. and foreign patents, maskwork rights,
//copyrights and other intellectual property laws.
//
//This reference design file, and your use thereof, is subject to and
//governed by the terms and conditions of the applicable Altera Reference
//Design License Agreement.  By using this reference design file, you
//indicate your acceptance of such terms and conditions between you and
//Altera Corporation.  In the event that you do not agree with such terms and
//conditions, you may not use the reference design file. Please promptly
//destroy any copies you have made.
//
//This reference design file being provided on an "as-is" basis and as an
//accommodation and therefore all warranties, representations or guarantees
//of any kind (whether express, implied or statutory) including, without
//limitation, warranties of merchantability, non-infringement, or fitness for
//a particular purpose, are specifically disclaimed.  By making this
//reference design file available, Altera expressly does not recommend,
//suggest or require that this reference design file be used in combination
//with any other product not provided by Altera
//----------------------------------------------------------------------------*/

//Group Enable Definitions
//This lists every pinout group
//Users can enable any group by uncommenting the corresponding line below:
//`define enable_ADC
//`define enable_ARDUINO
//`define enable_GPIO0
//`define enable_GPIO1
//`define enable_HPS

module fpga_main(
	//////////// CLOCK //////////
	input						FPGA_CLK_50,
	input						FPGA_CLK2_50,
	input						FPGA_CLK3_50,

`ifdef enable_ADC
	//////////// ADC //////////
	/* 3.3-V LVTTL */
	output						ADC_CONVST,
	output						ADC_SCLK,
	output						ADC_SDI,
	input						ADC_SDO,
`endif

`ifdef enable_ARDUINO
	//////////// ARDUINO ////////////
	/* 3.3-V LVTTL */
	inout					[15:0]	ARDUINO_IO,
	inout								ARDUINO_RESET_N,
`endif

`ifdef enable_GPIO0
	//////////// GPIO 0 ////////////
	/* 3.3-V LVTTL */
	inout				[35:0]		GPIO_0,
`endif

`ifdef enable_GPIO1
	//////////// GPIO 1 ////////////
	/* 3.3-V LVTTL */
	inout				[35:0]		GPIO_1,
`endif

`ifdef enable_HPS
	//////////// HPS //////////
	/* 3.3-V LVTTL */
	inout						HPS_CONV_USB_N,

	/* SSTL-15 Class I */
	output			[14:0]		HPS_DDR3_ADDR,
	output			 [2:0]		HPS_DDR3_BA,
	output						HPS_DDR3_CAS_N,
	output						HPS_DDR3_CKE,
	output						HPS_DDR3_CS_N,
	output			 [3:0]		HPS_DDR3_DM,
	inout			[31:0]		HPS_DDR3_DQ,
	output						HPS_DDR3_ODT,
	output						HPS_DDR3_RAS_N,
	output						HPS_DDR3_RESET_N,
	input						HPS_DDR3_RZQ,
	output						HPS_DDR3_WE_N,
	/* DIFFERENTIAL 1.5-V SSTL CLASS I */
	output						HPS_DDR3_CK_N,
	output						HPS_DDR3_CK_P,
	inout			 [3:0]		HPS_DDR3_DQS_N,
	inout			 [3:0]		HPS_DDR3_DQS_P,

	/* 3.3-V LVTTL */
	output						HPS_ENET_GTX_CLK,
	inout						HPS_ENET_INT_N,
	output						HPS_ENET_MDC,
	inout						HPS_ENET_MDIO,
	input						HPS_ENET_RX_CLK,
	input			 [3:0]		HPS_ENET_RX_DATA,
	input						HPS_ENET_RX_DV,
	output			 [3:0]		HPS_ENET_TX_DATA,
	output						HPS_ENET_TX_EN,
	inout						HPS_GSENSOR_INT,
	inout						HPS_I2C0_SCLK,
	inout						HPS_I2C0_SDAT,
	inout						HPS_I2C1_SCLK,
	inout						HPS_I2C1_SDAT,
	inout						HPS_KEY,
	inout						HPS_LED,
	inout						HPS_LTC_GPIO,
	output						HPS_SD_CLK,
	inout						HPS_SD_CMD,
	inout			 [3:0]		HPS_SD_DATA,
	output						HPS_SPIM_CLK,
	input						HPS_SPIM_MISO,
	output						HPS_SPIM_MOSI,
	inout						HPS_SPIM_SS,
	input						HPS_UART_RX,
	output						HPS_UART_TX,
	input						HPS_USB_CLKOUT,
	inout			 [7:0]		HPS_USB_DATA,
	input						HPS_USB_DIR,
	input						HPS_USB_NXT,
	output						HPS_USB_STP,
`endif

	//////////// KEY ////////////
	/* 3.3-V LVTTL */
	input				[1:0]			KEY,

	//////////// LED ////////////
	/* 3.3-V LVTTL */
	output				[7:0]			LED,

	//////////// SW ////////////
	/* 3.3-V LVTTL */
	input				[3:0]			SW

	/////////// USER ///////////

);

	assign LED[1:0] = SW[3:0];

	// assign ARR[0][0] = 1;
	// assign ARR[1][1] = 0;
	// assign ARR[2][2] = 1;

	// assign ARR[0][0] = (SW [0] && SW [1]);
	// assign ARR[0][1] = (SW [1] && SW [2]);
	// assign ARR[0][2] = (SW [2] && SW [3]);
	//
	// assign ARR[1][0] = (ARR[0][0] && ARR[0][1]);
	// assign ARR[1][1] = (ARR[0][1] && ARR[0][2]);
	//
	// assign ARR[2][0] = (ARR[1][0] && ARR[1][1]);
	//
	// assign LED [0]	= ARR[2][0];

endmodule
